module my100Hz (input logic clk, reset,
              output logic clk100Hz
             );
    logic q0,q1,q2,q3,q4,q5,q6,q7,q8,q9,q10,q11,q12,q13,q14,q15,q16;
    
    tflipflop ff0(
        .reset(reset),
        .clk(clk),
        .clk_out(q0)
    );
    tflipflop ff1(
        .reset(reset),
        .clk(q0),
        .clk_out(q1)
    );
    tflipflop ff2(
        .reset(reset),
        .clk(q1),
        .clk_out(q2)
    );
    tflipflop ff3(
        .reset(reset),
        .clk(q2),
        .clk_out(q3)
    );
    tflipflop ff4(
        .reset(reset),
        .clk(q3),
        .clk_out(q4)
    );
    tflipflop ff5(
        .reset(reset),
        .clk(q4),
        .clk_out(q5)
    );
    tflipflop ff6(
        .reset(reset),
        .clk(q5),
        .clk_out(q6)
    );
    tflipflop ff7(
        .reset(reset),
        .clk(q6),
        .clk_out(q7)
    );
    tflipflop ff8(
        .reset(reset),
        .clk(q7),
        .clk_out(q8)
    );
    tflipflop ff9(
        .reset(reset),
        .clk(q8),
        .clk_out(q9)
    );
    tflipflop ff10(
        .reset(reset),
        .clk(q9),
        .clk_out(q10)
    );
    tflipflop ff11(
        .reset(reset),
        .clk(q10),
        .clk_out(q11)
    );
    tflipflop ff12(
        .reset(reset),
        .clk(q11),
        .clk_out(q12)
    );
    tflipflop ff13(
        .reset(reset),
        .clk(q12),
        .clk_out(q13)
    );
    tflipflop ff14(
        .reset(reset),
        .clk(q13),
        .clk_out(q14)
    );
    tflipflop ff15(
        .reset(reset),
        .clk(q14),
        .clk_out(q15)
    );
    tflipflop ff16(
        .reset(reset),
        .clk(q15),
        .clk_out(q16)
    );
    tflipflop ff17(
        .reset(reset),
        .clk(q16),
        .clk_out(q17)
    );
    tflipflop ff18(
        .reset(reset),
        .clk(q17),
        .clk_out(q18)
    );
    tflipflop ff19(
        .reset(reset),
        .clk(q18),
        .clk_out(clk100Hz)
    );

endmodule